`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/06/19 14:24:40
// Design Name: 
// Module Name: and_gate
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//------------------------------------------------------------------------------------------------------------//
module and_gate(
    input A,
    input B,
    output F
    );
    
    and(F, A, B);    //��ȣ�� �� ó���� ���   and���� �⺻���� ���� �����Ǿ� ����  and(a,b,c)�� ���� ���� ���� ������ �ʰ� �׳� ����ϸ� ��
    
endmodule 
//------------------------------------------------------------------------------------------------------------//
module half_adder_structural(    //structural("������ �𵨸�")   half_adder(�ݰ����) sum = 2�Է� ���� ��� carry  = 2�Է� ������ �� �߻��ϴ� �ø� ��
    input A,                     
    input B,
    output sum,                       //00 - 0  /   01 - 1  /  10   -  1   / 11 - 0
    output carry                       //00 - 0  /  01 - 0    / 10   -  0  /  11 - 1
    );
    
    xor(sum, A, B);
    and(carry, A, B);
    
endmodule
//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module half_adder(    //dataflow modeling(�����Ͱ� ��� �귯������ ���)
    input A,
    input B,
    output sum,
    output carry
    );
    
    assign sum = A ^ B;         //^ = XOR   assign�� ����ϸ� ������ �÷ο� �𵨸���
    assign carry = A & B;       //& = AND
    
endmodule
//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
//module h_adder(    
//        input A,
//        input B,
//        output sum,
//        output carry
//);

//        assign sum = ({A,B} == 2'b00) ? 0 : ({A,B} == 2'b11) ? 0 : 1;
//        assign carry = ({A,B} == 2'b11) ? 1 : 0;
        
//endmodule
//------------------------------------------------------------------------------------------------------------//
module half_adder_behavioral(    //  "������ �𵨸�" ->�߻��� ǥ��
    input A,
    input B,
    output reg sum,             // reg : ��������Type���� �ٲ��ִ� �Լ�
    output reg carry
    );
    
    always @(A, B)begin
        case({A, B})                                                    //��� �Է¿� ���ؼ� �� �����ؾ��� or default�� ����ϸ� ��(�������� ���� ������ ���� default�� ��)
            2'b00: begin sum = 0; carry = 0; end           //gate�� ������ �����ϴ� �� (������ �𵨸�)
            2'b01: begin sum = 1; carry = 0; end           //������ ������ ��������Type�̾����
            2'b10: begin sum = 1; carry = 0; end           //��Ʈ ���� ������ ���� ������ 2'b �� ���� 2��Ʈ ���̳ʸ��� ���� ǥ����
            2'b11: begin sum = 0; carry = 1; end           // {} : ���տ����ڷ� ��� // C����� {}�� verilog������ begin - end�� ǥ����
                                                                                    //MUX�� ������
        endcase
    end
endmodule
//------------------------------------------------------------------------------------------------------------//
//������� ����� ������ ����Ʈ�� ����� ���� "�ν��Ͻ�ȭ"
//�������� �ݰ���⸦ 2�� �����
module full_adder_structural(                 //������ �𵨸����� ������ �� ������ �𵨸� ���X
    input A, B, cin,
    output sum, carry
    );
    
    wire sum_0, carry_0;            //half_adder�� sum, carry ����� ��Ÿ�� ����
    wire carry_1;
    
    half_adder ha0 (.A(A), .B(B), .sum(sum_0), .carry(carry_0));          //�ν��Ͻ��� ���鶧 .A��� �ϸ� "half_adder"�� ����� ������ ����
                                                                                                                            //(A) ��ȣ���� A�� ���� "full_adder"�� ����� ������ ����
                                                                                                                 //�����ϸ� half_adder�� A�� full_adder�� A�� �״�� ��(B�� ��������)
    half_adder ha1 (.A(sum_0), .B(cin), .sum(sum), .carry(carry_1));
                                                                                                                    //.A(sum_0) -> half_adder�� A�� full_adder�� sum_0������ �������� ���� ����
    
    or (carry, carry_0, carry_1);
endmodule
//------------------------------------------------------------------------------------------------------------//
//------------------------------------------------------------------------------------------------------------//
module f_add(       //4bit ������� ������ �÷ο� �𵨸�
        input [3:0] A, B,
        input C,
        output [3:0] sum,
        output carry 
);
        wire [4:0] temp;
        
        assign temp = A+B+C;
        assign sum = temp[3:0];
        assign carry = temp[4];

endmodule
//------------------------------------------------------------------------------------------------------------//
module f_add_top();
        reg [3:0] A, B;
        reg C;
        wire [3:0] sum;
        wire carry;
        
        

endmodule
//------------------------------------------------------------------------------------------------------------//
module full_adder(                 //������ �𵨸����� ������ ��
    input A, B, cin,
    output sum, carry
    );
    
    assign sum = A ^ B ^ cin;                                                                           //�Ϲ����� ���α׷� ���� ������ ���� ���۵��� ����
    assign carry = (cin & (A ^ B)) | (A & B);        //cin(A xor B) + AB      // ���ı����� ���ôٹ������� �����
    
    
endmodule
//------------------------------------------------------------------------------------------------------------//

//4bits ���İ���� : ������� 4���� ���ķ� ������ ȸ��  ripple carry adder(RCA)��� ��(carry�� �ѱ�� ���)
module fadder_4bit_structural(
    input [3:0] a, b,                 //0,1,2,3 bit�� ������ a�� �������   [�ֻ��� ��Ʈ(MSB) : ������ ��Ʈ(LSB)]
    input cin,
    output [3:0] sum,
    output carry
    );
    
    wire [2:0] carry_in;
    
    full_adder fa0 (.A(a[0]), .B(b[0]), .cin(cin), .sum(sum[0]), .carry(carry_in[0]));    
    full_adder fa1 (.A(a[1]), .B(b[1]), .cin(carry_in[0]), .sum(sum[1]), .carry(carry_in[1]));
    full_adder fa2 (.A(a[2]), .B(b[2]), .cin(carry_in[1]), .sum(sum[2]), .carry(carry_in[2]));
    full_adder fa3 (.A(a[3]), .B(b[3]), .cin(carry_in[2]), .sum(sum[3]), .carry(carry));
    
endmodule
//------------------------------------------------------------------------------------------------------------//
module fadder_4bit(         //������ �𵨸� full_adder
    input [3:0] a, b,                 //0,1,2,3 bit�� ������ a�� �������   [�ֻ��� ��Ʈ(MSB) : ������ ��Ʈ(LSB)]
    input cin,
    output [3:0] sum,
    output carry
    );
    
    wire [4:0] temp;
    
    assign temp = a + b + cin;          //4bit + 4bit + carry = 5bit
    assign sum = temp[3:0];            //���� 4��Ʈ�� sum
    assign carry = temp[4];              //�ֻ��� 1��Ʈ�� carry �� �ȴ�
    
endmodule
//------------------------------------------------------------------------------------------------------------//

//8��Ʈ �� �� �ֻ��� ��Ʈ�� 1�̸�(1000 0000 = -128(����)) �ֻ�����Ʈ�� 0�̸�(0111 1111 = 127(���)) 
// -> -128~127
//-1�� ǥ���� ���� -1�� ����� 1�� ��Ʈ���� ��Ų �� +1 ���ָ� ��
//-> 1000 0000(-1)�� ����� 0000 0001(1)�� ���� ��Ű�� 1111 1110 ���⿡ +1 = 1111 1111 -> 
//bit clear : AND, bit set : OR , bit toglle : XOR
//------------------------------------------------------------------------------------------------------------//
module fadd_sub_4bit_s(
    input [3:0] a, b,                 //0,1,2,3 bit�� ������ a�� �������   [�ֻ��� ��Ʈ(MSB) : ������ ��Ʈ(LSB)]
    input s,                                //s = 0(�����) , s = 1(�����)
    output [3:0] sum,
    output carry
    );
    
    wire [2:0] carry_in;
    
    full_adder fa0 (.A(a[0]), .B(b[0] ^ s), .cin(s), .sum(sum[0]), .carry(carry_in[0]));             //b�Է��� s�� XOR��
    full_adder fa1 (.A(a[1]), .B(b[1] ^ s), .cin(carry_in[0]), .sum(sum[1]), .carry(carry_in[1]));
    full_adder fa2 (.A(a[2]), .B(b[2] ^ s), .cin(carry_in[1]), .sum(sum[2]), .carry(carry_in[2]));
    full_adder fa3 (.A(a[3]), .B(b[3] ^ s), .cin(carry_in[2]), .sum(sum[3]), .carry(carry));
    
    
endmodule
//------------------------------------------------------------------------------------------------------------//

//SYNTHESIS : RTL(VHDL, Verilog source)�� gate level�� netlist�� ��ȯ�ϴ� �ܰ��Դϴ�.
//  �� ���� ������ RTL ���踦 power, timing�� ���� constraint�� ����Ͽ�
//     gate�� �̷���� netlist�� �ٲ��ִ� �߿��� �۾��Դϴ�.

//PDT ����Ʈ���� ���������ð��� ���� 
//�ִ뵿�����ļ��� �������� ����

//���ճ�ȸ�� : �Է¿� ���� ����� ������
//������ȸ�� : ���� ������ ��¿� ���� ����� ������(CLK�� ���)

//------------------------------------------------------------------------------------------------------------//
module fadd_sub_4bit(
    input [3:0] a, b,                 //0,1,2,3 bit�� ������ a�� �������   [�ֻ��� ��Ʈ(MSB) : ������ ��Ʈ(LSB)]
    input s,                                //s = 0(�����) , s = 1(�����)
    output [3:0] sum,
    output carry
    );
    
    wire [4:0] temp;                                     //5��Ʈ ¥��
    
    assign temp = s ? a - b:  a + b;                        //���ϱ��� ���     ���ǿ����� ?���� ���̸� : ������ temp�� ?���� �����̸� : �������� temp�� ��                       
    assign sum = temp[3:0];
    assign carry = temp[4];
    
    //���� ���� �˰�����
    
endmodule
//------------------------------------------------------------------------------------------------------------//


//------------------------------------------------------------------------------------------------------------//
module comparator (
            input A, B,
            output equal, greater, less
        );
        
    assign equal = A ~^ B;                  //assign���� ��������� �������𵨸��� ����
    assign greater = A & ~B;
    assign less = ~A & B;
    
endmodule
//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module comparator2 #(parameter N = 4)(              //N�� 4�� �ٲ�� compile ����
            input [N-1:0] A, B,
            output equal, greater, less
        );
        
    assign equal = (A == B) ? 1'b1 : 1'b0;                  //? : ���� ������ ���̸� : ���� 
    assign greater = (A > B) ? 1'b1 : 1'b0;
    assign less = (A < B)? 1'b1 : 1'b0;
    
endmodule
//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module decoder_2_4 (            
            input [1:0] A,
            output [3:0] Y

            );
            //������ �÷ο� �𵨸�
            assign Y = (A == 2'b00) ? 4'b0001 : (A == 2'b01) ? 4'b0010 : (A == 2'b10) ? 4'b0100 : 4'b1000;
            //?�� ���̸� ���� ���� �����̸� : �������� ���ǹ��� �߰��Ͽ� ��� �̾�� �� ����
            
            //���ڴ� ������ �𵨸�
//            always @(A) begin    //@(A) �� A�� �Է��� ���� --> always���� @(������ ������ ���� ���ϸ� �ѹ� �����Ѵ�)
//                    case(A)                 
//                        2'b00: Y = 4'b0001;     //A=00�̸�
//                        2'b01: Y = 4'b0010; 
//                        2'b10: Y = 4'b0100; 
//                        2'b11: Y = 4'b1000;
//                                                                        //���� A�� 4���� ���θ� ������� ������ ������ default���� ����� �����                                                
//                    endcase  
//            end

//            always @(A) begin    //@(A) �� A�� �Է��� ���� --> always���� @(������ ������ ���� ���ϸ� �ѹ� �����Ѵ�)
//                    if(A == 2'b00) Y = 4'b0001;
//                    else if(A == 2'b01) Y = 4'b0010;
//                    else if(A == 2'b10) Y = 4'b0100;
//                    else Y = 4'b1000;
//            end

endmodule
//------------------------------------------------------------------------------------------------------------//



//------------------------------------------------------------------------------------------------------------//

module decoder_2_4_en (            
            input [1:0] A,
            input en,
            output reg [3:0] Y

            );
            //������ �÷ο� �𵨸�
            //assign Y = (en == 0) ? 4'b0000 : (A == 2'b00) ? 4'b0001 : (A == 2'b01) ? 4'b0010 : (A == 2'b10) ? 4'b0100 : 4'b1000;
            //?�� ���̸� ���� ���� �����̸� : �������� ���ǹ��� �߰��Ͽ� ��� �̾�� �� ����
            
//            always @(A) begin    //@(A) �� A�� �Է��� ���� --> always���� @(������ ������ ���� ���ϸ� �ѹ� �����Ѵ�)
//                if(en == 1) begin
//                    case(A)                 
//                        2'b00: Y = 4'b0001;     //A=00�̸�
//                        2'b01: Y = 4'b0010; 
//                        2'b10: Y = 4'b0100; 
//                        2'b11: Y = 4'b1000;
//                                                                        //���� A�� 4���� ���θ� ������� ������ ������ default���� ����� �����                                                
//                    endcase  
//            end
//            else Y = 0;
//            end

            always @(A) begin    //@(A) �� A�� �Է��� ���� --> always���� @(������ ������ ���� ���ϸ� �ѹ� �����Ѵ�)
                if(en == 1)begin
                    if(A == 2'b00) Y = 4'b0001;
                    else if(A == 2'b01) Y = 4'b0010;
                    else if(A == 2'b10) Y = 4'b0100;
                    else Y = 4'b1000;
                end
                else Y = 0;
            end
            
endmodule

//------------------------------------------------------------------------------------------------------------//
module decoder_3_8 (                    //������ �𵨸����� 3X8���ڴ� ����
        input [2:0] D,
        output [7:0] Y
                
        );

        decoder_2_4_en de0 (.A(D[1:0]), .en(!D[2]), .Y(Y[3:0]));
        
        decoder_2_4_en de1 (.A(D[1:0]), .en(D[2]), .Y(Y[7:4]));

endmodule
//------------------------------------------------------------------------------------------------------------//


//------------------------------------------------------------------------------------------------------------//
module decoder_7seg(
                input [3:0] hex_value ,
                output reg [7:0] seg_7
);
                //������ �𵨸�
        always @(hex_value) begin
                case(hex_value)
                    4'b0000 : seg_7 = 8'b0000_0011;              //����ǥ�� A�� �ֻ�����Ʈ�� ���
                    4'b0001 : seg_7 = 8'b1001_1111;         //1
                    4'b0010 : seg_7 = 8'b0010_0101;         //2
                    4'b0011 : seg_7 = 8'b0000_1101;         //3
                    4'b0100 : seg_7 = 8'b1001_1001;         //4
                    4'b0101 : seg_7 = 8'b0100_1001;         //5
                    4'b0110 : seg_7 = 8'b0100_0001;         //6
                    4'b0111 : seg_7 = 8'b0001_1111;         //7
                    4'b1000 : seg_7 = 8'b0000_0001;         //8
                    4'b1001 : seg_7 = 8'b0000_1001;         //9
                    4'b1010 : seg_7 = 8'b0001_0001;         //A
                    4'b1011 : seg_7 = 8'b1100_0001;         //B
                    4'b1100 : seg_7 = 8'b0110_0011;         //C
                    4'b1101 : seg_7 = 8'b1000_0101;         //D
                    4'b1110 : seg_7 = 8'b0110_0001;         //E
                    4'b1111 : seg_7 = 8'b0111_0001;         //F
                    
                endcase
        end  

endmodule

//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module fnd_test_top(            //������ ����°� �������ִ� ��� : TOP
        input clk,                        //clk�� �ִٴ� ���� ������ȸ�ζ�� ����            
        output [7:0] seg_7,
        output [3:0] com        //4��Ʈ ¥�� FND�̹Ƿ� COM ���� 4�� �ʿ�
);
        
        assign com = 4'b0011;
        
        reg [25:0] clk_div;
        
        always @(posedge clk) clk_div = clk_div + 1;        //rising edge���� 26��Ʈ¥�� clk_div(reg)�� 1�� ���� ��Ų�� ���ֺ�
                                                                                    
        reg [3:0] count;
        always @(negedge clk_div[25])begin          //8ns X 2^26 ~= 0.5s
                count = count + 1;
        end
        //wire [7:0] seg_7_font;        common
    decoder_7seg seg7(.hex_value(count), .seg_7(seg_7));            //
        //assign seg_7 = ~seg_7_font;
endmodule
//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module encoder_4_2(           
            input [3:0] D,
            output [1:0] B
);

        assign B = (D == 4'b0001) ? 2'b00 : (D == 4'b0010) ? 2'b01 : (D == 4'b0100) ? 2'b10 : 2'b11;
        //���ڴ��� �Է��� �������ٴ� ���� �Ͽ� ����Ǿ���� ���⼭�� D�� 4�Է� �ܿ��� ���ٶ�� ������ �� ����
        //������ vivado ���α׷������� �Է��� 4���ۿ� ���´ٴ� ���� �𸣴� ������    -> �Է����� ������ ���� �ƴ� D���� ��� ���ǹ��� �� ���� 11�� ������

endmodule

//------------------------------------------------------------------------------------------------------------//


//------------------------------------------------------------------------------------------------------------//
module mux_2_1(
            input [1:0] d,
            input s,
            output f
);
            
            assign f = s ? d[1] : d[0];
endmodule
//������ �𵨸�
//        wire sbar, in0, in1;        
        
//        not (sbar, s);
//        and (in0, d[0], sbar);
//        and (in1, d[1], s);
//        or (f, in0, in1);


//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module mux_4_1(
            input [3:0] d,
            input [1:0] s,
            output f
);
            //assign f = s ? d[1] : d[0];
            //�����ϰ� �� �� ����
            assign f = d[s];        //�̷���               

endmodule


//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module mux_8_1(
            input [7:0] d,
            input [2:0] s,
            output f
);
            assign f = d[s];        //�̷���   s�� 3��Ʈ�� ��

endmodule


//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module demux_1_4(
        input d,
        input [1:0] s,
        output [3:0] f
//        output reg [3:0] f
);

//        always @*begin  //d�� s�� �ٲ�� always�� 1�� ����  always @(d, s)begin = always @*begin   * : �Է��� �����̶� ���ϸ� always�� 1�� ����
//            f = 0;              //f�� ������������ �κ��� 0���� ��
//            f[s] = d;       //s=0�̸� d�� f[0]���� s=1�̸� d�� f[1]�� ������ 
//        end

        assign f = (s == 2'b00) ? {3'b000, d} : (s == 2'b01) ? {2'b00, d, 1'b0} : (s == 2'b10) ? {1'b0, d, 2'b00} : {d, 3'b000};
endmodule
//------------------------------------------------------------------------------------------------------------//

//------------------------------------------------------------------------------------------------------------//
module mux_test_top(
        input [7:0] d,
        input [2:0] s_mux,
        input [1:0] s_demux,
        output [3:0] f
);

         wire w;                //mux�� ��� wire�ϳ� �ʿ�
         
         mux_8_1 mux(.d(d), .s(s_mux), .f(w));
       
         demux_1_4 demux(.d(w), .s(s_demux), .f(f));
        
        
endmodule
//------------------------------------------------------------------------------------------------------------//



































